`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:14:04 03/11/2015 
// Design Name: 
// Module Name:    mux2to1_32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mux2to1_32(input [31:0] a,
					  input [31:0] b,
					  input sel,
					  output [31:0] o
    );
	 
	 assign o = ({32{!sel}} & a) | ({32{sel}} & b);


endmodule
